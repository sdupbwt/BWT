`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07.05.2020 01:26:58
// Design Name: 
// Module Name: sort4elem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sort4elem(
//    input wire clk,
//    input wire rst,
//    input wire [7:0] array_L [INPUT_ARR_LEN-1:0],
//    input wire [7:0] array_R [INPUT_ARR_LEN-1:0],
//    output reg [7:0] [2*INPUT_ARR_LEN-1:0] merged_array 
    );
    
    
    
endmodule
